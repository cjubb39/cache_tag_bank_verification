bind l2_cache_tag_unisim_rtl l2_cache_tag_checker_sva check_1
(clk, rst, tag_in_valid, set_in_valid, 
state_in_valid, inv_ack_cnt_in_valid, 
flush_in_valid, flush_complete_ready, 
way_out_ready, state_out_ready, inv_ack_cnt_out_ready, tag_out_evict_ready, 
set_out_evict_ready, state_out_evict_ready, way_out_flush_ready, 
inv_ack_cnt_out_flush_ready, tag_out_flush_ready, set_out_flush_ready, 
state_out_flush_ready, 
internal_state,
tag_in_ready, set_in_ready, state_in_ready, 
inv_ack_cnt_in_ready, flush_in_ready, flush_complete_valid,
way_out_valid, state_out_valid,
inv_ack_cnt_out_valid, tag_out_evict_valid, 
set_out_evict_valid,
state_out_evict_valid, way_out_flush_valid, 
inv_ack_cnt_out_flush_valid,
tag_out_flush_valid, set_out_flush_valid,
state_out_flush_valid, mem_tag_CE0,
mem_tag_WE0, mem_tag_CE1, mem_tag_CE2, mem_tag_CE3, 
mem_tag_CE4, mem_tag_CE5, mem_tag_CE6, 
mem_tag_CE7, mem_tag_CE8, mem_state_CE0, 
mem_state_WE0, mem_state_CE1,
mem_state_CE2, mem_state_CE3, mem_state_CE4, 
mem_state_CE5, mem_state_CE6,
mem_state_CE7, mem_state_CE8, mem_inv_ack_cnt_CE0, 
mem_inv_ack_cnt_WE0, mem_inv_ack_cnt_CE1, 
mem_inv_ack_cnt_CE2, mem_inv_ack_cnt_CE3, 
mem_inv_ack_cnt_CE4, mem_inv_ack_cnt_CE5, 
mem_inv_ack_cnt_CE6, mem_inv_ack_cnt_CE7, 
mem_inv_ack_cnt_CE8);
